module exec_unit(
    input [1:0] databus_opcode,
    input [3:0] databus_addr,
    input [7:0] databus_datain,
    input [2:0] ALU_opcode,
    output [7:0] databus_dataout,
);
endmodule